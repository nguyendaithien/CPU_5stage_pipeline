`include "defi.vh"
module CPU_EDABK_TOP #( parameter DATA_WIDTH = 32) (
   clk
  ,rst_n
  ,RD
  ,WR
  ,A_DMEM
  ,A_IMEM // address
  ,Instr_in
  ,D_in
  ,D_out
  ,DMEM_rst
  ,byte_mark
  ,boot_add
 );

   input              clk       ;
   input              rst_n     ;
   output             RD        ;
   output             WR        ;
   input       [31:0] boot_add  ;
   input       [31:0] Instr_in  ;
   input       [31:0] D_in      ;
   output wire [31:0] A_DMEM    ;
   output wire [31:0] A_IMEM    ;
   output wire [31:0] D_out     ;
   output wire [2:0 ] byte_mark ;
   output wire        DMEM_rst  ;

 
   wire [4:0 ] WB_rd_add         ;
   wire [31:0] WB_data_write_reg ;
   wire        WB_regwrite       ;
   // output of IF stage
   wire [31:0] IF_instr          ;
   wire [4:0 ] IMEM_add          ;
   wire [31:0] IF_pc             ;
   // OUTPUT ID stage
   wire [4:0 ] ID_rs1_add        ;
   wire [4:0 ] ID_rs2_add        ;
   wire [4:0 ] ID_rd_add         ;
   wire [31:0] ID_rs1_data       ;
   wire [31:0] ID_rs2_data       ;
   wire [31:0] ID_pc             ;
   wire [3:0 ] ID_alu_op         ;
   wire [31:0] ID_imm            ;
   wire [1:0 ] ID_sel_to_reg     ;
   wire        ID_regwrite       ;
   wire [3:0 ] mem_op            ;
   wire        ID_jump           ;
   wire ID_RD                    ;
   wire ID_WR                    ;
   wire        ID_branch         ;
   wire [1:0 ] ID_alu_sel1       ;
   wire [1:0 ] ID_alu_sel2       ;
   wire        ID_pc_sel         ;
   // OUTPUT EX stage
   wire [31:0] EX_pc             ;
   wire [4:0 ] EX_rs1_add        ;
   wire [4:0 ] EX_rs2_add        ;
   wire [4:0 ] EX_rd_add         ;
   wire [1:0 ] EX_sel_to_reg     ;
   wire        EX_regwrite       ;
   wire        EX_RD             ;
   wire        EX_WR             ;
   wire [3:0 ] EX_mem_op         ;
   wire [31:0] EX_alu_result     ;
   wire        EX_zero           ;
   wire [31:0] EX_imm            ;
   wire [31:0] EX_pc_dest        ;
   wire [31:0] EX_rs2_data       ;
   // output of MEM stage
   wire [31:0] MEM_add           ;
   wire [3:0 ] DMEM_byte_mark    ;
   wire [31:0] DMEM_data_write   ;
   wire [31:0] MEM_data          ;
   wire        MEM_regwrite      ;
   wire [31:0] MEM_alu_result    ;
   wire [4:0 ] MEM_rd_add        ;
   wire [1:0 ] MEM_sel_to_reg    ;
   wire        MEM_RD_mem        ;
   wire        MEM_WR_mem        ;
   wire [31:0] MEM_pc            ;

  IF_stage #( .DATA_WIDTH(32))  if_stage (
     .clk        (clk         )
    ,.rst_n      (rst_n       )
    ,.IF_instr_i (            )
    ,.boot_add   (boot_add    )
    ,.flush      (IF_ID_flush )
    ,.pc_dest    (EX_pc_dest  )
    ,.IMEM_data_i(Instr_in    )
    ,.stall      (stall       )
    ,.pc_sel     (ID_pc_sel   )
    ,.IF_pc_o    (IF_pc       )
    ,.IF_instr_o (IF_instr    )
    ,.IMEM_add_o (A_IMEM      )
  );


  ID_stage #( .DATA_WIDTH(32)) id_stage (
   .clk            (clk           ) 
  ,.rst_n          (rst_n         )
  ,.stall          (stall         )
  ,.flush          (IF_ID_flush   )
  ,.ID_instr_i     (IF_instr      )
  ,.EX_ALU_result_i(EX_alu_result )
  ,.EX_rd_add_i    (EX_rd_add     )
  ,.WB_data_i      (WB_data       )
  ,.WB_regwrite_i  (WB_regwrite   )
  ,.WB_rd_add_i    ( WB_rd_add    )
  ,.ID_pc_i        (IF_pc         )
  ,.ID_rs1_add_o   (ID_rs1_add    )
  ,.ID_rs2_add_o   (ID_rs2_add    )
  ,.ID_rd_add_o    (ID_rd_add     )
  ,.ID_rs1_data_o  (ID_rs1_data   )
  ,.ID_rs2_data_o  (ID_rs2_data   )
  ,.ID_pc_o        (ID_pc         )
  ,.ID_imm_o       (ID_imm        )
  ,.ID_alu_op_o    (ID_alu_op     )
  ,.ID_regwrite_o  (ID_regwrite   )
  ,.ID_mem_op_o    (ID_mem_op     )
  ,.ID_jump_o      (ID_jump       )
  ,.ID_sel_to_reg_o(ID_sel_to_reg )
  ,.ID_RD_en_o     (ID_RD         )
  ,.ID_WR_en_o     (ID_WR         )
  ,.ID_branch_o    (ID_branch     )
  ,.ID_alu_sel1_o  (ID_alu_sel1   )
  ,.ID_alu_sel2_o  (ID_alu_sel2   )
  ,.ID_pc_sel_o    (ID_pc_sel     )
);


  EX_stage #( .DATA_WIDTH(32)) ex_stage (
     .clk             (clk               )                               
    ,.rst_n           (rst_n             )
    ,.EX_pc_i         (ID_pc             )
    ,.EX_rs1_add_i    (ID_rs1_add        )
    ,.EX_rs2_add_i    (ID_rs2_add        )
    ,.EX_rd_add_i     (ID_rd_add         )
    ,.EX_sel_to_reg_i (ID_sel_to_reg     )
    ,.EX_regwrite_i   (ID_regwrite       )
    ,.EX_RD_mem_i     (ID_RD             )
    ,.EX_WR_mem_i     (ID_WR             )
    ,.EX_mem_op_i     (ID_mem_op         )
    ,.EX_rs2_data_i   (ID_rs2_data       )
    ,.EX_rs1_data_i   (ID_rs1_data       )
    ,.EX_sel_alu1_i   (EX_alu_sel1       )
    ,.EX_sel_alu2_i   (EX_alu_sel2       )
    ,.EX_imm_i        (ID_imm            )
    ,.flush           (EX_flush          )
    ,.forwardA        (forward_A         )
    ,.forwardB        (forward_B         )
    ,.WB_data_i       (WB_data_write_reg )
    ,.EX_data_i       (EX_alu_result     )
    ,.hazard          (                  )
    ,.EX_rs2_data_o   (EX_rs2_data       )
    ,.EX_pc_o         (EX_pc             )
    ,.EX_rs1_add_o    (EX_rs1_add        )
    ,.EX_rs2_add_o    (EX_rs2_add        )
    ,.EX_rd_add_o     (EX_rd_add         )
    ,.EX_sel_to_reg_o (EX_sel_to_reg     )
    ,.EX_regwrite_o   (EX_regwrite       )
    ,.EX_RD_mem_o     (EX_RD             )
    ,.EX_WR_mem_o     (EX_WR             )
    ,.EX_mem_op_o     (EX_mem_op         )
    ,.EX_alu_result_o (EX_alu_result     )
    ,.EX_zero_o       (EX_zero           )
    ,.EX_imm_o        (EX_imm            )
    ,.EX_pc_dest      (EX_pc_dest        )
);

   MEM_stage #( .DATA_WIDTH(32)) mem_stage (
     .clk               (clk               )
    ,.rst_n             (rst_n             )
    ,.WB_data_i         (WB_data_write_reg )
    ,.forward           (                  )
    ,.MEM_RD_mem_i      (EX_RD             )
    ,.MEM_WR_mem_i      (EX_WR             )
    ,.MEM_mem_op_i      (EX_mem_op         )
    ,.MEM_regwrite_i    (EX_regwrite       )
    ,.MEM_alu_result_i  (EX_alu_result     )
    ,.MEM_rs2_data_i    (EX_rs2_data       )
    ,.MEM_rd_add_i      (EX_rd_add         )
    ,.MEM_pc_i          (EX_pc             )
    ,.MEM_imm_i         (EX_imm            )
    ,.MEM_imm_o         (MEM_imm           )
    ,.MEM_pc_o          (MEM_pc            )
    ,.DMEM_add_o        (M_add             )
    ,.DMEM_byte_mark_o  (DMEM_byte_mark    )
    ,.DMEM_data_write_o (DMEM_data_write   )
    ,.MEM_data_o        (MEM_data          )
    ,.MEM_regwrite_o    (MEM_regwrite      )
    ,.MEM_alu_result_o  (MEM_alu_result    )
    ,.MEM_rd_add_o      (MEM_rd_add        )
    ,.MEM_sel_to_reg_o  (MEM_sel_to_reg    )
    ,.MEM_sel_to_reg_i  (EX_sel_to_reg     )
    ,.MEM_RD_mem_o      (MEM_RD_mem        )
    ,.MEM_WR_mem_o      (MEM_WR_mem        )
    ,.DMEM_data_i       (D_in              ) // data from DMEM
    ,.DMEM_rst_o        (DMEM_rst          )
  );

  WB_stage #(.DATA_WIDTH(32))  wb_stage (
   .clk                   (clk               )
  ,.rst_n                 (rst_n             )
  ,.WB_rd_add_i           (MEM_rd_add        )
  ,.DMEM_data_i           (MEM_data          )
  ,.WB_alu_result_i       (MEM_alu_result    )
  ,.WB_sel_to_reg_i       (MEM_sel_to_reg    )
  ,.WB_regwrite_i         (MEM_regwrite      )
  ,.WB_pc_i               (MEM_pc            )
  ,.WB_imm_i              (MEM_imm           )
  ,.WB_rd_add_o           (WB_rd_add         )
  ,.WB_data_write_reg_o   (WB_data_write_reg )
  ,.WB_regwrite_o         (WB_regwrite       )
  );


   CONTROL_HAZARD #( .DATA_WIDTH(32)) control_hazard (
   .clk(clk)
  ,.rst_n          (rst_n        )
  ,.stall_o        (stall        )
  ,.IF_ID_flush_o  (IF_ID_flush  )
  ,.EX_flush_o     (EX_flush     )
  ,.hazard         (hazard       )
  ,.forward_A_o    (forward_A    )
  ,.forward_B_o    (forward_B    )
  ,.forward_dmem   (forward_dmem )
  ,.ID_RD_mem_i    (ID_RD        )
  ,.ID_rs1_add_i   (ID_rs1_add   )
  ,.ID_rs2_add_i   (ID_rs2_add   )
  ,.ID_rd_add_i    (ID_rd_add    )
  ,.EX_rs1_add_i   (EX_rs1_add   )
  ,.EX_rs2_add_i   (EX_rs2_add   )
  ,.EX_rd_add_i    (EX_rd_add    )
  ,.MEM_rd_add_i   (MEM_rd_add   )
  ,.EX_regwrite_i  (EX_regwrite  )
  ,.MEM_regwrite_i (MEM_regwrite )
  ,.IF_instr_i     (IF_instr     )
  ,.ID_jump        (ID_jump      )
  ,.zero           (EX_zero      )
 );

 endmodule



