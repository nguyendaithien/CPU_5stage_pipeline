coverpoint mode {
 bins zero = {0}; 
 bins zero = {1}; 

 bins range[] = {[0:$]};

 bins c[] = {[2:3] , [5,7] };

 bins range[4] = { [0:$]};

 bins range[4] = { [],1,3,6 };

 bins orthers = default;
}
  
  
